library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_signed.all;
entity button is
  port (
    pSW0 : IN std_logic;
    pSW1 : IN std_logic;
    pSW2 : IN std_logic;
    pSW3 : IN std_logic
  );
end button;

architecture RTL of button is

begin  -- RTL

  

end RTL;
